module main;
  initial
    begin
      $display("Howdy Hackers");
      $finish;
    end
endmodule
